* NGSPICE file created from addf.ext - technology: sky130A

.subckt addf A S CO vdd gnd B CI
X0 a_952_521# CI a_870_521# vdd sky130_fd_pr__pfet_01v8 ad=0.164 pd=1.52 as=0.164 ps=1.52 w=1.26 l=0.15
X1 S a_784_115# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.334 pd=3.05 as=0.214 ps=1.6 w=1.26 l=0.15
X2 a_526_115# CI gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X3 a_27_521# B vdd vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X4 a_952_115# CI a_870_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0676 pd=0.78 as=0.0676 ps=0.78 w=0.52 l=0.15
X5 S a_784_115# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.57 as=0.0884 ps=0.86 w=0.52 l=0.15
X6 vdd A a_27_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.334 ps=3.05 w=1.26 l=0.15
X7 a_784_115# CON a_526_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X8 a_27_115# B gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X9 gnd A a_27_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.138 ps=1.57 w=0.52 l=0.15
X10 a_784_115# CON a_526_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X11 CON CI a_27_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X12 vdd A a_368_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.132 ps=1.47 w=1.26 l=0.15
X13 a_526_521# A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X14 CO CON vdd vdd sky130_fd_pr__pfet_01v8 ad=0.334 pd=3.05 as=0.334 ps=3.05 w=1.26 l=0.15
X15 CON CI a_27_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X16 a_870_521# B a_784_115# vdd sky130_fd_pr__pfet_01v8 ad=0.164 pd=1.52 as=0.176 ps=1.54 w=1.26 l=0.15
X17 gnd A a_368_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0546 ps=0.73 w=0.52 l=0.15
X18 a_526_115# A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X19 CO CON gnd gnd sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.57 as=0.138 ps=1.57 w=0.52 l=0.15
X20 a_870_115# B a_784_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0676 pd=0.78 as=0.0728 ps=0.8 w=0.52 l=0.15
X21 a_368_521# B CON vdd sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.47 as=0.176 ps=1.54 w=1.26 l=0.15
X22 vdd B a_526_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X23 vdd A a_952_521# vdd sky130_fd_pr__pfet_01v8 ad=0.214 pd=1.6 as=0.164 ps=1.52 w=1.26 l=0.15
X24 a_368_115# B CON gnd sky130_fd_pr__nfet_01v8 ad=0.0546 pd=0.73 as=0.0728 ps=0.8 w=0.52 l=0.15
X25 gnd B a_526_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X26 gnd A a_952_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0884 pd=0.86 as=0.0676 ps=0.78 w=0.52 l=0.15
X27 a_526_521# CI vdd vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
C0 CON a_368_115# 0.0037f
C1 a_526_115# a_368_115# 6.28e-19
C2 CON a_526_115# 0.0428f
C3 CON a_27_521# 0.066f
C4 vdd a_952_521# 0.00964f
C5 a_784_115# a_526_521# 0.0546f
C6 CON a_27_115# 0.0441f
C7 CON a_368_521# 0.00367f
C8 a_27_115# a_27_521# 0.00483f
C9 a_784_115# vdd 0.149f
C10 S B 8.48e-19
C11 CON a_952_115# 0.00227f
C12 a_784_115# a_870_521# 0.0133f
C13 S A 0.0302f
C14 a_526_521# CI 0.023f
C15 CO S 0.0234f
C16 a_784_115# a_870_115# 0.00424f
C17 vdd CI 0.122f
C18 CI a_870_521# 0.00263f
C19 a_784_115# CON 0.169f
C20 a_784_115# a_526_115# 0.0359f
C21 a_526_521# B 0.036f
C22 a_784_115# a_368_521# 5.73e-19
C23 vdd B 0.293f
C24 a_526_521# A 0.00216f
C25 CON CI 0.216f
C26 a_784_115# a_952_115# 0.00282f
C27 a_870_521# B 0.0013f
C28 a_526_115# CI 0.0258f
C29 a_27_521# CI 0.00307f
C30 vdd A 0.167f
C31 vdd CO 0.112f
C32 a_27_115# CI 0.00565f
C33 a_870_115# B 2.05e-19
C34 a_784_115# a_952_521# 0.0127f
C35 CI a_952_115# 5.65e-19
C36 a_368_115# B 9.37e-19
C37 CON B 0.281f
C38 a_526_115# B 0.0263f
C39 a_27_521# B 0.0591f
C40 CON A 0.453f
C41 a_952_521# CI 0.00174f
C42 a_526_521# S 6.86e-19
C43 CON CO 0.127f
C44 a_27_115# B 0.0277f
C45 a_368_521# B 0.00709f
C46 a_526_115# A 0.00873f
C47 a_27_521# A 0.0145f
C48 vdd S 0.14f
C49 a_27_115# A 0.0428f
C50 a_784_115# CI 0.0932f
C51 S a_870_521# 7.59e-19
C52 a_952_115# A 3.88e-19
C53 S a_870_115# 3.84e-19
C54 a_952_521# A 0.00141f
C55 CON S 0.113f
C56 a_784_115# B 0.19f
C57 a_27_521# S 2.01e-19
C58 a_526_521# vdd 0.175f
C59 a_784_115# A 0.19f
C60 S a_368_521# 1.28e-19
C61 a_784_115# CO 0.00108f
C62 CI B 0.879f
C63 S a_952_115# 7.1e-19
C64 vdd a_870_521# 0.0066f
C65 CI A 0.533f
C66 CO CI 4.26e-19
C67 a_526_521# CON 0.00605f
C68 a_952_521# S 0.00114f
C69 a_526_521# a_526_115# 0.00723f
C70 vdd a_368_115# 1.02e-19
C71 CON vdd 0.17f
C72 a_784_115# S 0.116f
C73 vdd a_526_115# 0.00164f
C74 a_27_521# vdd 0.133f
C75 A B 0.513f
C76 a_27_115# vdd 8.57e-19
C77 vdd a_368_521# 0.00893f
C78 CO B 0.00429f
C79 CON a_870_115# 0.00202f
C80 S CI 0.00855f
C81 CO A 6.94e-19
.ends

